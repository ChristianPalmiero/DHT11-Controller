library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity dht11_sa is
  generic(
    freq:    positive range 1 to 1000 -- Clock frequency (MHz)
  );
  port(
    clk:      in  std_ulogic;
    rst:      in  std_ulogic;                    -- Active high synchronous reset
    btn:      in  std_ulogic;
    sw:       in  std_ulogic_vector(3 downto 0); -- Slide switches
    data_in:  in  std_ulogic;
    data_drv: out std_ulogic;
    led:      out std_ulogic_vector(3 downto 0)  -- LEDs
  );
end entity dht11_sa;

architecture rtl of dht11_sa is

  signal start             : std_ulogic;
  signal pe                : std_ulogic;
  signal b		   : std_ulogic;
  signal do                : std_ulogic_vector(39 downto 0);
  signal sipo_out_mux_in   : std_ulogic_vector(31 downto 0);
  signal checksum          : std_ulogic_vector(7 downto 0);
  signal checksum_ver_to_B : std_ulogic_vector(3 downto 0);
  signal nib_sel_to_A      : std_ulogic_vector(3 downto 0);

begin

  deb: entity work.debouncer(rtl)
  port map(
    clk   => clk,
    rst   => rst,
    d     => btn,
    q     => open,
    r     => start,
    f     => open,
    a     => open
  );

  u0: entity work.dht11_ctrl(rtl)
  generic map(
    freq => freq
  )
  port map(
    clk      => clk,
    srstn    => NOT(rst),
    start    => start,
    data_in  => data_in,
    data_drv => data_drv,
    pe       => pe,
    b        => b,
    do       => do
  );

  sipo_out_mux_in <= do(39 DOWNTO 8);
  checksum <= do(7 DOWNTO 0);

  MUXes: process(sipo_out_mux_in, sw)
  begin
    nib_sel_to_A <= sipo_out_mux_in(3 DOWNTO 0) when SW(0)='0' and SW(1)='0' and SW(2)='0' else
    sipo_out_mux_in(7 DOWNTO 4) when SW(0)='0' and SW(1)='0' and SW(2)='1' else
    sipo_out_mux_in(11 DOWNTO 8) when SW(0)='0' and SW(1)='1' and SW(2)='0' else
    sipo_out_mux_in(15 DOWNTO 12) when SW(0)='0' and SW(1)='1' and SW(2)='1' else
    sipo_out_mux_in(19 DOWNTO 16) when SW(0)='1' and SW(1)='0' and SW(2)='0' else
    sipo_out_mux_in(23 DOWNTO 20) when SW(0)='1' and SW(1)='0' and SW(2)='1' else
    sipo_out_mux_in(27 DOWNTO 24) when SW(0)='1' and SW(1)='1' and SW(2)='0' else
    sipo_out_mux_in(31 DOWNTO 28) when SW(0)='1' and SW(1)='1' and SW(2)='1';
  end process MUXes;

  Checksum_controller: process(checksum, sipo_out_mux_in)
  variable sum: std_ulogic_vector(7 DOWNTO 0);
  begin
    sum:= sipo_out_mux_in(31 DOWNTO 24) + sipo_out_mux_in(23 DOWNTO 16) + sipo_out_mux_in(15 DOWNTO 8) + sipo_out_mux_in(7 DOWNTO 0);
    if sum = checksum then
      checksum_ver_to_B(0) <= '0';
    else
      checksum_ver_to_B(0) <= '1';
    end if;
  end process Checksum_controller;

  checksum_ver_to_B(1) <= b;
  checksum_ver_to_B(2) <= SW(0);
  checksum_ver_to_B(3) <= pe;

  MUX: process(nib_sel_to_A, checksum_ver_to_B, SW(3))
  begin
    led <= nib_sel_to_A when (SW(3) = '1') else checksum_ver_to_B;
  end process MUX;

end architecture rtl;
